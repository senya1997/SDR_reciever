module fifo_async(

);



endmodule 
